//QR_Engine FSM
`define init        0
`define load_h      1
`define load_y      2
`define last_trig   3

//cal_Rii module FSM
`define idle 	    0
`define cal_sum     1
`define cal_sqrt    2
`define root1       1
`define root2       2
//y_process module FSM
`define idle 	    0
`define mult_QY_1   1
`define mult_QY_2   2

`define expan_bit   10   
